
module lab7_soc (
	clk_clk,
	game_rst_sig,
	key_external_connection_export,
	keycode_export,
	led_wire_export,
	leds_export,
	move_ready,
	move_hl_export,
	reset_reset_n,
	reset_game_export,
	reset_sw_export,
	sdram_clk_clk,
	sdram_wire_addr,
	sdram_wire_ba,
	sdram_wire_cas_n,
	sdram_wire_cke,
	sdram_wire_cs_n,
	sdram_wire_dq,
	sdram_wire_dqm,
	sdram_wire_ras_n,
	sdram_wire_we_n,
	spi0_MISO,
	spi0_MOSI,
	spi0_SCLK,
	spi0_SS_n,
	start_sw_export,
	text_ctrl_keycode,
	usb_gpx_export,
	usb_irq_export,
	usb_rst_export,
	vga_port_blue,
	vga_port_green,
	vga_port_red,
	vga_port_hs,
	vga_port_vs,
	win_export,
	win_cond_edge,
	menu_hex,
	sw_digits_export);	

	input		clk_clk;
	output		game_rst_sig;
	input	[1:0]	key_external_connection_export;
	output	[7:0]	keycode_export;
	output	[7:0]	led_wire_export;
	output	[13:0]	leds_export;
	input		move_ready;
	output		move_hl_export;
	input		reset_reset_n;
	input		reset_game_export;
	output		reset_sw_export;
	output		sdram_clk_clk;
	output	[12:0]	sdram_wire_addr;
	output	[1:0]	sdram_wire_ba;
	output		sdram_wire_cas_n;
	output		sdram_wire_cke;
	output		sdram_wire_cs_n;
	inout	[15:0]	sdram_wire_dq;
	output	[1:0]	sdram_wire_dqm;
	output		sdram_wire_ras_n;
	output		sdram_wire_we_n;
	input		spi0_MISO;
	output		spi0_MOSI;
	output		spi0_SCLK;
	output		spi0_SS_n;
	output		start_sw_export;
	input	[7:0]	text_ctrl_keycode;
	input		usb_gpx_export;
	input		usb_irq_export;
	output		usb_rst_export;
	output	[3:0]	vga_port_blue;
	output	[3:0]	vga_port_green;
	output	[3:0]	vga_port_red;
	output		vga_port_hs;
	output		vga_port_vs;
	output		win_export;
	input		win_cond_edge;
	output	[3:0]	menu_hex;
	input	[15:0]	sw_digits_export;
endmodule
